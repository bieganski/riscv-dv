/home/mateusz/github/mtkcpu/mtkcpu/tests/riscv_dv_assets/riscv_core_setting.sv